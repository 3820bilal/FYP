module tb_upcounter (
input	logic			clk,
input	logic			reset,

);
endmodule