module Baseboard (
input	logic		clk,
input	logic		reset

);
endmodule