module clock (
input	logic		clk,
input	logic		reset,
output	logic	[5:0]	count_sec,
output	logic	[5:0]	count_min,
output	logic	[5:0]	count_hrs

);
endmodule