module AND
(
	input	a,
	input	b,
	output reg c
);

always@*
c = a & b;

endmodule