module test (
input	logic		clk,
input	logic		reset,
input	logic		inp1
);

endmodule