module Baseboard (
input	logic			clk,
input	logic			reset,

);


counter bilal
(
.clk			(),
.reset			(),
.en			(),
.clr			(),
.count			()
);

endmodule